library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
--use IEEE.NUMERIC_STD.ALL;

entity bit_cntr is
--  Port ( );
end bit_cntr;

architecture arch of bit_cntr is

begin


end arch;