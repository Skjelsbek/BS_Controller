library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
--use IEEE.NUMERIC_STD.ALL;

entity deserializer is
--  Port ( );
end deserializer;

architecture arch of deserializer is

begin


end arch;
