library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
--use IEEE.NUMERIC_STD.ALL;

entity prog_cntr is
--  Port ( );
end prog_cntr;

architecture arch of prog_cntr is

begin


end arch;