library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
--use IEEE.NUMERIC_STD.ALL;

entity latch is
--  Port ( );
end latch;

architecture arch of latch is

begin


end arch;