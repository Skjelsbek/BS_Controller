library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
--use IEEE.NUMERIC_STD.ALL;

entity fsm is
--  Port ( );
end fsm;

architecture arch of fsm is

begin


end arch;
