library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
--use IEEE.NUMERIC_STD.ALL;

entity shift_cntr is
--  Port ( );
end shift_cntr;

architecture arch of shift_cntr is

begin


end arch;