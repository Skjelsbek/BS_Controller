library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
--use IEEE.NUMERIC_STD.ALL;

entity ins_reg_tb is
--  Port ( );
end ins_reg_tb;

architecture arch of ins_reg_tb is

begin


end arch;