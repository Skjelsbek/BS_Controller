library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
--use IEEE.NUMERIC_STD.ALL;

entity comparator_tb is
--  Port ( );
end comparator_tb;

architecture arch of comparator_tb is

begin

end arch;