library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
--use IEEE.NUMERIC_STD.ALL;

entity fsm_tb is
--  Port ( );
end fsm_tb;

architecture arch of fsm_tb is

begin


end arch;