library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
--use IEEE.NUMERIC_STD.ALL;

entity comparator is
--  Port ( );
end comparator;

architecture arch of comparator is

begin


end arch;