library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
--use IEEE.NUMERIC_STD.ALL;

entity bs_controller_tb is
--  Port ( );
end bs_controller_tb;

architecture arch of bs_controller_tb is

begin


end arch;
