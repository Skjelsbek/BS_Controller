library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
--use IEEE.NUMERIC_STD.ALL;

entity prog_cntr_tb is
--  Port ( );
end prog_cntr_tb;

architecture arch of prog_cntr_tb is

begin


end arch;