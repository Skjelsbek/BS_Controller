library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
--use IEEE.NUMERIC_STD.ALL;

entity serializer_tb is
--  Port ( );
end serializer_tb;

architecture arch of serializer_tb is

begin


end arch;