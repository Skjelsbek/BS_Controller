library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
--use IEEE.NUMERIC_STD.ALL;

entity shift_cntr_tb is
--  Port ( );
end shift_cntr_tb;

architecture arch of shift_cntr_tb is

begin


end arch;