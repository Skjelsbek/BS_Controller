library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
--use IEEE.NUMERIC_STD.ALL;

entity serializer is
--  Port ( );
end serializer;

architecture arch of serializer is

begin


end arch;