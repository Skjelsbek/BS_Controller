library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
--use IEEE.NUMERIC_STD.ALL;

entity ins_reg is
--  Port ( );
end ins_reg;

architecture arch of ins_reg is

begin


end arch;