library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
--use IEEE.NUMERIC_STD.ALL;

entity latch_tb is
--  Port ( );
end latch_tb;

architecture arch of latch_tb is

begin


end arch;